library verilog;
use verilog.vl_types.all;
entity \_xor\ is
    port(
        result          : out    vl_logic;
        input1          : in     vl_logic;
        input2          : in     vl_logic
    );
end \_xor\;
