library verilog;
use verilog.vl_types.all;
entity MIPS_32bit_testbench is
end MIPS_32bit_testbench;
