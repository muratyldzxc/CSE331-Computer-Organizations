library verilog;
use verilog.vl_types.all;
entity MIPS_32bit is
    port(
        clock           : in     vl_logic
    );
end MIPS_32bit;
